package cache_types;

typedef logic [127:0] cache_line;
typedef logic [8:0] cache_tag;
typedef logic [2:0] cache_index;
typedef logic [3:0] cache_offset;
typedef logic [2:0] cache_read_offset;

endpackage : cache_types